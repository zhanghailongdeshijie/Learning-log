`timescale       1ns/1ns

module  tb_clk_gen();

reg     sys_clk     ;
reg     sys_rst_n   ;
wire     inclk0      ;
wire     areset      ;

wire    c0          ;
wire    locked      ;


initial
    begin
        sys_clk = 1'b1;
        sys_rst_n <= 1'b0;
        #20
        sys_rst_n <= 1'b1;
    end
    
always #10 sys_clk = ~sys_clk;

clk_gen     tb_clk_gen_
(
    .sys_clk        (sys_clk  ),
    .sys_rst_n      (sys_rst_n),

    .inclk0         (inclk0   ),
    .areset         (areset   ),

    .c0             (c0       ),
    .locked         (locked   )

);

endmodule